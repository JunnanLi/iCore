/*
 *  TuMan32 -- A Small but pipelined RISC-V (RV32I) Processor Core
 *  Copyright (C) 2019-2020 Junnan Li <lijunnan@nudt.edu.cn>
 *
 *  Permission to use, copy, modify, and/or distribute this code for any purpose with or
 *   without fee is hereby granted, provided that the above copyright notice and this 
 *   permission notice appear in all copies.
 *
 *	Function description: This module is used to generate FAST packets to configure itcm 
 *	 and dtcm of CPU.
 */
`timescale 1 ns / 1 ps

module gen_data(
	input 					clk,
	input 					resetn,

	output	reg 			data_in_valid,
	output	reg 	[133:0]	data_in,
	input					data_out_valid,
	input			[133:0]	data_out
);
	/** regs:
	*		memory[64KB] used to store instruction; 
	*/
	
	wire [1023:0][31:0] memory = {
		32'h0040006f,
		32'h00000093,
		32'h00000113,
		32'h00000193,
		32'h00000213,
		32'h00000293,
		32'h00000313,
		32'h00000393,
		32'h00000413,
		32'h00000493,
		32'h00000513,
		32'h00000593,
		32'h00000613,
		32'h00000693,
		32'h00000713,
		32'h00000793,
		32'h00000813,
		32'h00000893,
		32'h00000913,
		32'h00000993,
		32'h00000a13,
		32'h00000a93,
		32'h00000b13,
		32'h00000b93,
		32'h00000c13,
		32'h00000c93,
		32'h00000d13,
		32'h00000d93,
		32'h00000e13,
		32'h00000e93,
		32'h00000f13,
		32'h00000f93,
		32'h00010137,
		32'hdeadc1b7,
		32'heef18193,
		32'h00018213,
		32'h044000ef,
		32'h10000537,
		32'h04400593,
		32'h04f00613,
		32'h04e00693,
		32'h04500713,
		32'h00a00793,
		32'h00b52023,
		32'h00c52023,
		32'h00d52023,
		32'h00e52023,
		32'h00f52023,
		32'h20000537,
		32'h075bd5b7,
		32'hd1558593,
		32'h00b52023,
		32'h00100073,
		32'hff010113,
		32'h2c800513,
		32'h00112623,
		32'h048000ef,
		32'h00001737,
		32'h800066b7,
		32'h80000637,
		32'h00100593,
		32'h00300513,
		32'h80070713,
		32'h00c68693,
		32'h00c60793,
		32'h0007a803,
		32'h00b81463,
		32'h00a7a023,
		32'h00e787b3,
		32'hfed798e3,
		32'hfe9ff06f,
		32'h100007b7,
		32'h00a7a023,
		32'h00008067,
		32'h10000737,
		32'h00054783,
		32'h00079463,
		32'h00008067,
		32'h00150513,
		32'h00f72023,
		32'hfedff06f,
		32'hfe010113,
		32'h00812c23,
		32'h00410413,
		32'h00912a23,
		32'h01212823,
		32'h00112e23,
		32'h00050493,
		32'h00040913,
		32'h02049c63,
		32'h03240a63,
		32'h10000737,
		32'hfff44783,
		32'hfff40413,
		32'h03078793,
		32'h00f72023,
		32'hff2418e3,
		32'h01c12083,
		32'h01812403,
		32'h01412483,
		32'h01012903,
		32'h02010113,
		32'h00008067,
		32'h00a00593,
		32'h00048513,
		32'h0a4000ef,
		32'h00a40023,
		32'h00a00593,
		32'h00048513,
		32'h04c000ef,
		32'h00140413,
		32'h00050493,
		32'hfa5ff06f,
		32'hfff58593,
		32'h00259593,
		32'h2f800713,
		32'h100006b7,
		32'h0005d463,
		32'h00008067,
		32'h00b557b3,
		32'h00f7f793,
		32'h00f707b3,
		32'h0007c783,
		32'hffc58593,
		32'h00f6a023,
		32'hfe1ff06f,
		32'h06054063,
		32'h0605c663,
		32'h00058613,
		32'h00050593,
		32'hfff00513,
		32'h02060c63,
		32'h00100693,
		32'h00b67a63,
		32'h00c05863,
		32'h00161613,
		32'h00169693,
		32'hfeb66ae3,
		32'h00000513,
		32'h00c5e663,
		32'h40c585b3,
		32'h00d56533,
		32'h0016d693,
		32'h00165613,
		32'hfe0696e3,
		32'h00008067,
		32'h00008293,
		32'hfb5ff0ef,
		32'h00058513,
		32'h00028067,
		32'h40a00533,
		32'h0005d863,
		32'h40b005b3,
		32'hf9dff06f,
		32'h40b005b3,
		32'h00008293,
		32'hf91ff0ef,
		32'h40a00533,
		32'h00028067,
		32'h00008293,
		32'h0005ca63,
		32'h00054c63,
		32'hf79ff0ef,
		32'h00058513,
		32'h00028067,
		32'h40b005b3,
		32'hfe0558e3,
		32'h40a00533,
		32'hf61ff0ef,
		32'h40b00533,
		32'h00028067,
		32'h00001941,
		32'h73697200,
		32'h01007663,
		32'h0000000f,
		32'h33767205,
		32'h70326932,
		32'h00000030,
		32'h4347000a,
		32'h28203a43,
		32'h29554e47,
		32'h322e3920,
		32'h4100302e,
		32'h0000001b,
		32'h63736972,
		32'h11010076,
		32'h04000000,
		32'h76720510,
		32'h32693233,
		32'h00003070,
		32'h33323130,
		32'h37363534,
		32'h42413938,
		32'h46454443,
		32'h00000000,
		32'h00001b41,
		32'h73697200,
		32'h01007663,
		32'h00000011,
		32'h72051004,
		32'h69323376,
		32'h00307032,
		32'h00001941,
		32'h73697200,
		32'h01007663,
		32'h0000000f,
		32'h33767205,
		32'h70326932,
		32'h00000030,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0
    };

	// reg 	[31:0] 	memory [0:64*1024/4-1];
	
	reg 	[13:0] 	addr_q;
    wire 	[31:0]	memory_data;
    reg 	[31:0]	addr_conf;

    reg 	[3:0]	count,pkt_count;

     always @* begin
    	addr_q <= 13'h3ff - addr_conf[9:0];
    end
	assign memory_data = memory[addr_q];

	reg [4:0]	state_mem;
	parameter 	IDLE_S 		= 5'd0,
				FAKE_DATA_S	= 5'd1,
				CONF_TCM_S	= 5'd2,
				CONF_TCM_1_S= 5'd3,
				CONF_TCM_2_S= 5'd4,
				CONF_SEL_1_S= 5'd5,
				CONF_SEL_2_S= 5'd6,
				READY_S		= 5'd7,
				READ_1_S	= 5'd8,
				READ_2_S	= 5'd9,
				READ_3_S	= 5'd10,
				READ_4_S	= 5'd11,
				READ_5_S	= 5'd12,
				READ_6_S	= 5'd13,
				WRITE_END_S	= 5'd14,
				WAIT_10_CLK_S= 5'd15,
				TEST_L2SW_S	= 5'd16;

	always @(posedge clk or negedge resetn) begin
		if (!resetn) begin
			// reset
//			addr_q 		<= 14'h400;
			state_mem 	<= IDLE_S;

			data_in_valid	<= 1'b0;
			data_in 		<= 134'b0;
			count			<= 4'b0;
			pkt_count		<= 4'b0;
			addr_conf		<= 32'b0;
		end
		else begin
			case(state_mem)
				IDLE_S: begin
					data_in_valid 	<= 1'b1;
					data_in 		<= {2'b01,4'b0,128'b0};
					state_mem 		<= FAKE_DATA_S;
					count 			<= 4'b0;
				end
				FAKE_DATA_S: begin
					count <= count + 4'd1;
					case(count)
						4'd0: data_in <= {2'b11, 4'b0, 128'd0};
						4'd1: data_in <= {2'b11, 4'b0, 96'b0,16'h9001,16'b0};
						4'd2: data_in <= {2'b11, 4'b0, 112'd1,16'b0};
						4'd3: data_in <= {2'b11, 4'b0, 112'd2,16'b0};
						4'd4: data_in <= {2'b11, 4'b0, 112'd3,16'b0};
						4'd5: data_in <= {2'b10, 4'b0, 112'd4,16'b0};
						default: begin
						end
					endcase
					if(count == 4'd5)
						state_mem <= CONF_TCM_S;
				end
				CONF_TCM_S: begin
					data_in_valid 	<= 1'b1;
					data_in 		<= {2'b01,4'b0,128'b0};
					state_mem 		<= CONF_TCM_1_S;
					count 			<= 4'b0;
				end
				CONF_TCM_1_S: begin
					count <= count + 4'd1;
					case(count)
						4'd0: data_in <= {2'b11, 4'b0, 128'd0};
						4'd1: data_in <= {2'b11, 4'b0, 96'b0,16'h9003,16'b0};
						default: begin
						end
					endcase
					if(count == 4'd1)
						state_mem <= CONF_TCM_2_S;
					//addr_q <= 14'h3ff;
					addr_conf <= 32'b0;
				end
				CONF_TCM_2_S: begin
					addr_conf 	<= addr_conf + 32'd1;
					//addr_q 		<= addr_q - 14'd1;
					data_in[131:0] <= {4'b0, 48'd0, memory_data, addr_conf,16'b0};
					if(addr_conf == 32'd1023) begin
						state_mem <= READ_1_S;
						data_in[133:132] <= {2'b10};
					end
					else begin
						state_mem <= CONF_TCM_2_S;
						data_in[133:132] <= {2'b11};
					end
				end
				CONF_SEL_1_S: begin
					data_in_valid 	<= 1'b1;
					data_in 		<= {2'b01,4'b0,128'b0};
					state_mem 		<= CONF_SEL_2_S;
					count 			<= 4'b0;
				end
				CONF_SEL_2_S: begin
					count <= count + 4'd1;
					case(count)
						4'd0: data_in <= {2'b11, 4'b0, 128'd0};
						4'd1: data_in <= {2'b11, 4'b0, 96'b0,16'h9001,16'b0};
						4'd2: data_in <= {2'b11, 4'b0, 128'd0};
						4'd3: data_in <= {2'b11, 4'b0, 128'd1};
						4'd4: data_in <= {2'b11, 4'b0, 128'd2};
						4'd5: data_in <= {2'b10, 4'b0, 128'd3};
						default: begin
						end
					endcase
					if(count == 4'd5) begin
						count		<= 4'd0;
						state_mem 	<= WAIT_10_CLK_S;
					end
				end
				READ_1_S: begin
					data_in_valid 	<= 1'b1;
					data_in 		<= {2'b01,4'b0,128'b0};
					state_mem 		<= READ_2_S;
					count 			<= 4'b0;
				end
				READ_2_S: begin
					count <= count + 4'd1;
					case(count)
						4'd0: data_in <= {2'b11, 4'b0, 128'd0};
						4'd1: data_in <= {2'b11, 4'b0, 96'b0,16'h9002,16'b0};
						4'd2: data_in <= {2'b11, 4'b0, 128'd1};
						4'd3: data_in <= {2'b11, 4'b0, 128'd2};
						4'd4: data_in <= {2'b11, 4'b0, 128'd3};
						4'd5: data_in <= {2'b10, 4'b0, 128'd4};
						default: begin
						end
					endcase
					if(count == 4'd5)
						state_mem <= READ_3_S;
				end
				READ_3_S: begin
					data_in_valid 	<= 1'b1;
					data_in 		<= {2'b01,4'b0,128'b0};
					state_mem 		<= READ_4_S;
					count 			<= 4'b0;
				end
				READ_4_S: begin
					count <= count + 4'd1;
					case(count)
						4'd0: data_in <= {2'b11, 4'b0, 128'd0};
						4'd1: data_in <= {2'b11, 4'b0, 96'b0,16'h9004,16'b0};
						4'd2: data_in <= {2'b11, 4'b0, 112'd128,16'b0};
						4'd3: data_in <= {2'b11, 4'b0, 128'd2};
						4'd4: data_in <= {2'b11, 4'b0, 128'd3};
						4'd5: data_in <= {2'b10, 4'b0, 128'd4};
						default: begin
						end
					endcase
					if(count == 4'd5)
						state_mem <= READ_5_S;
				end
				READ_5_S: begin
					data_in_valid 	<= 1'b1;
					data_in 		<= {2'b01,4'b0,128'b0};
					state_mem 		<= READ_6_S;
					count 			<= 4'b0;
				end
				READ_6_S: begin
					count <= count + 4'd1;
					case(count)
						4'd0: data_in <= {2'b11, 4'b0, 128'd0};
						4'd1: data_in <= {2'b11, 4'b0, 96'b0,16'h9004,16'b0};
						4'd2: data_in <= {2'b11, 4'b0, 112'd129,16'b0};
						4'd3: data_in <= {2'b11, 4'b0, 128'd2};
						4'd4: data_in <= {2'b11, 4'b0, 128'd3};
						4'd5: data_in <= {2'b10, 4'b0, 128'd4};
						default: begin
						end
					endcase
					if(count == 4'd5)
						state_mem <= CONF_SEL_1_S;
				end
				WAIT_10_CLK_S: begin
					data_in_valid		<= 1'b0;
					count 				<= count + 4'd1;
					if(count == 4'd10) begin
						count 			<= 4'd0;
						data_in_valid 	<= 1'b1;
						data_in 		<= {2'b01,4'b0,128'b0};
						state_mem		<= TEST_L2SW_S;
					end
					else 
						state_mem		<= WAIT_10_CLK_S;
				end
				TEST_L2SW_S: begin
					count <= count + 4'd1;
					case(count)
						4'd0: data_in <= {2'b11, 4'b0, 128'd0};
						4'd1: data_in <= {2'b11, 4'b0, 96'b0,16'h0800,16'b0};
						4'd2: data_in <= {2'b11, 4'b0, 64'd6,64'd0};
						4'd3: data_in <= {2'b11, 4'b0, 128'd1};
						4'd4: data_in <= {2'b11, 4'b0, 128'd2};
						4'd5: data_in <= {2'b10, 4'b0, 128'd3};
						default: begin
						end
					endcase
					if(count == 4'd5) begin
						count			<= 4'd0;
						if(pkt_count == 4'd4)
							state_mem	<= READY_S;
						else begin
							state_mem 	<= WAIT_10_CLK_S;
							pkt_count	<= 4'd1 + pkt_count;
						end
					end
				end
				READY_S: begin
					data_in_valid <= 1'b0;
					state_mem <= READY_S;
				end
				default: begin
					state_mem <= IDLE_S;
				end
			endcase
		end
	end


endmodule