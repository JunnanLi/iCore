/*
 *  iCore_hardware -- Hardware for TuMan RISC-V (RV32I) Processor Core.
 *
 *  Copyright (C) 2019-2020 Junnan Li <lijunnan@nudt.edu.cn>.
 *  Copyright and related rights are licensed under the MIT license.
 *
 *	Data: 2020.01.01
 *	Description: This module is used to generate FAST packets to configure 
 *	 itcm and dtcm of CPU.
 *	Note: You can gen "gen_data_fixed_instr.sv" by running "write_instr.py"
 */
`timescale 1 ns / 1 ps


module gen_data(
	input 					clk,
	input 					resetn,

	output	reg 			data_in_valid,
	output	reg 	[133:0]	data_in,
	input					data_out_valid,
	input			[133:0]	data_out
);
	/** regs:
	*		memory[64KB] used to store instruction; 
	*/
	
	wire [2047:0][31:0] memory = {
		/**write_fix_instr*/
		32'h0040006f,
		32'h00000093,
		32'h00000113,
		32'h00000193,
		32'h00000213,
		32'h00000293,
		32'h00000313,
		32'h00000393,
		32'h00000413,
		32'h00000493,
		32'h00000513,
		32'h00000593,
		32'h00000613,
		32'h00000693,
		32'h00000713,
		32'h00000793,
		32'h00000813,
		32'h00000893,
		32'h00000913,
		32'h00000993,
		32'h00000a13,
		32'h00000a93,
		32'h00000b13,
		32'h00000b93,
		32'h00000c13,
		32'h00000c93,
		32'h00000d13,
		32'h00000d93,
		32'h00000e13,
		32'h00000e93,
		32'h00000f13,
		32'h00000f93,
		32'h00010137,
		32'hdeadc1b7,
		32'heef18193,
		32'h00018213,
		32'h044000ef,
		32'h10000537,
		32'h04400593,
		32'h04f00613,
		32'h04e00693,
		32'h04500713,
		32'h00a00793,
		32'h00b52023,
		32'h00c52023,
		32'h00d52023,
		32'h00e52023,
		32'h00f52023,
		32'h20000537,
		32'h075bd5b7,
		32'hd1558593,
		32'h00b52023,
		32'h00100073,
		32'h00002537,
		32'hf8010113,
		32'h89450513,
		32'h06112e23,
		32'h06812c23,
		32'h0c4000ef,
		32'h000017b7,
		32'h38978793,
		32'h00f11523,
		32'h0f82d7b7,
		32'hac578793,
		32'h04410513,
		32'h00000593,
		32'h00f12623,
		32'h679000ef,
		32'h00410593,
		32'h04410513,
		32'h6b1000ef,
		32'h000015b7,
		32'h01200613,
		32'h7d458593,
		32'h01c10513,
		32'h154000ef,
		32'h01600613,
		32'h00000593,
		32'h02e10513,
		32'h168000ef,
		32'h01c10593,
		32'h01400613,
		32'h04410513,
		32'h040010ef,
		32'h01c10593,
		32'h01400613,
		32'h04410513,
		32'h090010ef,
		32'h00050413,
		32'h00001537,
		32'h7bc50513,
		32'h040000ef,
		32'h07010793,
		32'h00878433,
		32'h01c10513,
		32'hfa040623,
		32'h02c000ef,
		32'h04410513,
		32'h0ec010ef,
		32'h14c000ef,
		32'h07c12083,
		32'h07812403,
		32'h08010113,
		32'h00008067,
		32'h100007b7,
		32'h00a7a023,
		32'h00008067,
		32'h10000737,
		32'h00054783,
		32'h00079463,
		32'h00008067,
		32'h00150513,
		32'h00f72023,
		32'hfedff06f,
		32'hfe010113,
		32'h00812c23,
		32'h00410413,
		32'h00912a23,
		32'h01212823,
		32'h00112e23,
		32'h00050493,
		32'h00040913,
		32'h02049c63,
		32'h03240a63,
		32'h10000737,
		32'hfff44783,
		32'hfff40413,
		32'h03078793,
		32'h00f72023,
		32'hff2418e3,
		32'h01c12083,
		32'h01812403,
		32'h01412483,
		32'h01012903,
		32'h02010113,
		32'h00008067,
		32'h00a00593,
		32'h00048513,
		32'h514010ef,
		32'h00a40023,
		32'h00a00593,
		32'h00048513,
		32'h4bc010ef,
		32'h00140413,
		32'h00050493,
		32'hfa5ff06f,
		32'hfff58593,
		32'h00002737,
		32'h00259593,
		32'h82c70713,
		32'h100006b7,
		32'h0005d463,
		32'h00008067,
		32'h00b557b3,
		32'h00f7f793,
		32'h00f707b3,
		32'h0007c783,
		32'hffc58593,
		32'h00f6a023,
		32'hfe1ff06f,
		32'h00000793,
		32'h00c79463,
		32'h00008067,
		32'h00f58733,
		32'h00074683,
		32'h00f50733,
		32'h00178793,
		32'h00d70023,
		32'hfe5ff06f,
		32'h00c50633,
		32'h00050793,
		32'h00c79463,
		32'h00008067,
		32'h00178793,
		32'hfeb78fa3,
		32'hff1ff06f,
		32'h200007b7,
		32'h0007a703,
		32'h00e52023,
		32'h0047a783,
		32'h00f52223,
		32'h00008067,
		32'h00002537,
		32'hff010113,
		32'h84050513,
		32'h00112623,
		32'hec5ff0ef,
		32'h00c12083,
		32'hf00007b7,
		32'h00100713,
		32'h00e7a023,
		32'h01010113,
		32'h00008067,
		32'hf9010113,
		32'h05512a23,
		32'h00058a93,
		32'h000025b7,
		32'h06812423,
		32'h06912223,
		32'h05612823,
		32'h00060493,
		32'h93458b13,
		32'h04000613,
		32'h93458593,
		32'h00050413,
		32'h01010513,
		32'h06112623,
		32'h07212023,
		32'h05312e23,
		32'h00078913,
		32'h00068993,
		32'h05412c23,
		32'h00070a13,
		32'hf2dff0ef,
		32'h01000613,
		32'h040b0593,
		32'h00010513,
		32'hf1dff0ef,
		32'h0024d603,
		32'h0044d783,
		32'h0009d503,
		32'h01061613,
		32'h00f66633,
		32'h0029d783,
		32'h00295803,
		32'h01051513,
		32'h00f56533,
		32'h00100793,
		32'h0004d883,
		32'h00095583,
		32'h01081813,
		32'h0cfa9063,
		32'hffff06b7,
		32'h00010737,
		32'h00d8e6b3,
		32'h00e8e733,
		32'h00d12a23,
		32'h00c12c23,
		32'h02e12223,
		32'h02c12423,
		32'h02a12623,
		32'h02b12a23,
		32'h80001737,
		32'h00241513,
		32'h82070713,
		32'h03012c23,
		32'h00e50733,
		32'h00000793,
		32'h04000693,
		32'h01010593,
		32'h00f585b3,
		32'h0005a583,
		32'h00f70633,
		32'h00478793,
		32'h00b62023,
		32'hfed794e3,
		32'h800017b7,
		32'h80078793,
		32'h00f50533,
		32'h01000713,
		32'h00000793,
		32'h00f10633,
		32'h00062603,
		32'h00f506b3,
		32'h00478793,
		32'h00c6a023,
		32'hfee796e3,
		32'h06812403,
		32'h06c12083,
		32'h06412483,
		32'h06012903,
		32'h05c12983,
		32'h05812a03,
		32'h05412a83,
		32'h05012b03,
		32'h00002537,
		32'h86850513,
		32'h07010113,
		32'hd55ff06f,
		32'h000a5683,
		32'h002a5783,
		32'h00c12c23,
		32'h01069693,
		32'h00f6e6b3,
		32'h004a5783,
		32'h00d12823,
		32'h02c12423,
		32'h01079793,
		32'h0117e733,
		32'h00e12a23,
		32'h00020737,
		32'h00e8e733,
		32'h00b7e7b3,
		32'h02e12223,
		32'h02a12623,
		32'h02d12823,
		32'h02f12a23,
		32'hf25ff06f,
		32'h00058793,
		32'h800005b7,
		32'h02e5d883,
		32'hfe010113,
		32'h00050713,
		32'h00001537,
		32'h00112e23,
		32'h00c12623,
		32'h80650513,
		32'h0aa89e63,
		32'h02c5d883,
		32'h00100313,
		32'hfff00513,
		32'h08689663,
		32'h0445de03,
		32'h0006d303,
		32'h086e1063,
		32'h04a5de03,
		32'h0026d303,
		32'h00d12423,
		32'h066e1863,
		32'h0245d503,
		32'h00a71023,
		32'h02a5d503,
		32'h00a71123,
		32'h0285d503,
		32'h00e12223,
		32'h00a71223,
		32'h03e5d503,
		32'h00a79023,
		32'h03c5d503,
		32'h00f12023,
		32'h00a79123,
		32'h00400513,
		32'h00a5a623,
		32'h0365d583,
		32'h03159e63,
		32'h00002537,
		32'h87450513,
		32'hc69ff0ef,
		32'h00012783,
		32'h00412703,
		32'h00812683,
		32'h00c12603,
		32'h00000513,
		32'h00200593,
		32'hda5ff0ef,
		32'h00100513,
		32'h01c12083,
		32'h02010113,
		32'h00008067,
		32'h00002537,
		32'h89850513,
		32'hc31ff0ef,
		32'h00200513,
		32'hfe5ff06f,
		32'hfff00513,
		32'hfddff06f,
		32'hf6010113,
		32'h09612023,
		32'h00002b37,
		32'h934b0b13,
		32'h08812c23,
		32'h08912a23,
		32'h09312623,
		32'h00050413,
		32'h00058993,
		32'h00060493,
		32'h050b0593,
		32'h07000613,
		32'h01010513,
		32'h08112e23,
		32'h09212823,
		32'h09412423,
		32'h09512223,
		32'h00070913,
		32'h00068a93,
		32'h00078a13,
		32'hca1ff0ef,
		32'h01000613,
		32'h0c0b0593,
		32'h00010513,
		32'h80098993,
		32'hc8dff0ef,
		32'h10099a63,
		32'h00095703,
		32'h00295783,
		32'h002a5503,
		32'h01071713,
		32'h00f76733,
		32'h00e12823,
		32'h00495703,
		32'h0004d783,
		32'h01051513,
		32'h01071713,
		32'h00f76733,
		32'h00e12a23,
		32'h0024d703,
		32'h0044d783,
		32'h00800593,
		32'h01071713,
		32'h00f76733,
		32'h000ad783,
		32'h00e12c23,
		32'h5a6c0737,
		32'h00e7e7b3,
		32'h002ad703,
		32'h02f12423,
		32'h000a5783,
		32'h01071713,
		32'h00f76733,
		32'h000017b7,
		32'h80078793,
		32'h00f56533,
		32'h02e12623,
		32'h02a12823,
		32'hbd1ff0ef,
		32'h80001737,
		32'h00241513,
		32'h82070713,
		32'h00e50733,
		32'h00000793,
		32'h07000693,
		32'h01010593,
		32'h00f585b3,
		32'h0005a583,
		32'h00f70633,
		32'h00478793,
		32'h00b62023,
		32'hfed794e3,
		32'h800017b7,
		32'h80078793,
		32'h00f50533,
		32'h01000713,
		32'h00000793,
		32'h00f10633,
		32'h00062603,
		32'h00f506b3,
		32'h00478793,
		32'h00c6a023,
		32'hfee796e3,
		32'h00002537,
		32'h8a850513,
		32'h09812403,
		32'h09c12083,
		32'h09412483,
		32'h09012903,
		32'h08c12983,
		32'h08812a03,
		32'h08412a83,
		32'h08012b03,
		32'h0a010113,
		32'haa5ff06f,
		32'h00002537,
		32'h8c450513,
		32'hfd1ff06f,
		32'h800006b7,
		32'h00050713,
		32'h0226d803,
		32'h00055503,
		32'h02068793,
		32'h06a81463,
		32'h0206d803,
		32'h00275683,
		32'hfff00513,
		32'h04d81e63,
		32'h0067d683,
		32'h00475703,
		32'h04e69863,
		32'h00e7d703,
		32'h80070713,
		32'h04071263,
		32'h0227d683,
		32'h0025d703,
		32'h02e69c63,
		32'h0267d683,
		32'h00065703,
		32'h02e69663,
		32'h0147c683,
		32'h00600713,
		32'h20000537,
		32'h00e69e63,
		32'h02c7d503,
		32'h100007b7,
		32'h01f57513,
		32'h00f50533,
		32'h00008067,
		32'hfff00513,
		32'h00008067,
		32'h00052703,
		32'h00100793,
		32'h0af71e63,
		32'hfe010113,
		32'h00912a23,
		32'h00050493,
		32'h00002537,
		32'h8e450513,
		32'h00812c23,
		32'h01212823,
		32'h00112e23,
		32'h01312623,
		32'h01448413,
		32'h9ddff0ef,
		32'h02448913,
		32'h00042503,
		32'h00800593,
		32'h00440413,
		32'ha65ff0ef,
		32'hff2418e3,
		32'h00002937,
		32'h89490513,
		32'h9b9ff0ef,
		32'h03448993,
		32'h00042503,
		32'h00800593,
		32'h00440413,
		32'ha41ff0ef,
		32'hff3418e3,
		32'h89490513,
		32'h999ff0ef,
		32'h04448913,
		32'h00042503,
		32'h00800593,
		32'h00440413,
		32'ha21ff0ef,
		32'hfe8918e3,
		32'h00002537,
		32'h8f450513,
		32'h975ff0ef,
		32'h01c12083,
		32'h01812403,
		32'h00400793,
		32'h00f4a023,
		32'h01012903,
		32'h01412483,
		32'h00c12983,
		32'h02010113,
		32'h00008067,
		32'h00008067,
		32'h800007b7,
		32'h00c7a683,
		32'h00100713,
		32'h00e69c63,
		32'h00300713,
		32'h00002537,
		32'h00e7a623,
		32'h90850513,
		32'h929ff06f,
		32'h00008067,
		32'h00000713,
		32'h00000793,
		32'h00b74e63,
		32'h0107d513,
		32'h00f50533,
		32'hfff54513,
		32'h01051513,
		32'h01055513,
		32'h00008067,
		32'h00171693,
		32'h00d506b3,
		32'h0006d683,
		32'h00170713,
		32'h00d787b3,
		32'hfd1ff06f,
		32'hfe010113,
		32'h00812c23,
		32'h80000437,
		32'h01512223,
		32'h00065703,
		32'h00068a93,
		32'h02245683,
		32'h00112e23,
		32'h00912a23,
		32'h01212823,
		32'h01312623,
		32'h01412423,
		32'h01612023,
		32'h1ae69263,
		32'h02045683,
		32'h00265703,
		32'h00050993,
		32'h00060913,
		32'hfff00513,
		32'h14e69863,
		32'h02645683,
		32'h00465703,
		32'h14e69263,
		32'h02e45703,
		32'h80070713,
		32'h12071c63,
		32'h03444683,
		32'h00100713,
		32'h12e69663,
		32'h02445703,
		32'h04045483,
		32'h03842b03,
		32'h00e99023,
		32'h02a45703,
		32'h00058a13,
		32'h00e99123,
		32'h02845703,
		32'h00e99223,
		32'h03845703,
		32'h00e59023,
		32'h03e45783,
		32'h00f59123,
		32'h80048793,
		32'h10079c63,
		32'h00002537,
		32'h91050513,
		32'h82dff0ef,
		32'h0009d783,
		32'h0029d703,
		32'hffff06b7,
		32'h01079793,
		32'h00e7e7b3,
		32'h02f42023,
		32'h0049d783,
		32'h00095703,
		32'h00db7b33,
		32'h01079793,
		32'h00e7e7b3,
		32'h02f42223,
		32'h00295783,
		32'h00495703,
		32'h01079793,
		32'h00e7e7b3,
		32'h000ad703,
		32'h02f42423,
		32'h002ad783,
		32'h01676733,
		32'h02e42c23,
		32'h000a5703,
		32'h01079793,
		32'h00e7e7b3,
		32'h002a5703,
		32'h02f42e23,
		32'h01071713,
		32'h04e42023,
		32'h03042583,
		32'h03042783,
		32'h0105d593,
		32'hfec58593,
		32'h0015d593,
		32'h0015f713,
		32'h02071063,
		32'h0107d793,
		32'hfec78793,
		32'hffc7f793,
		32'h00f40433,
		32'h04042783,
		32'h00d7f7b3,
		32'h04f42023,
		32'h80000437,
		32'h04442783,
		32'h04440513,
		32'h01079793,
		32'h0107d793,
		32'h04f42223,
		32'he49ff0ef,
		32'h04442783,
		32'h01051513,
		32'h00f56533,
		32'h04a42223,
		32'h00300793,
		32'h00f42623,
		32'h00048513,
		32'h01c12083,
		32'h01812403,
		32'h01412483,
		32'h01012903,
		32'h00c12983,
		32'h00812a03,
		32'h00412a83,
		32'h00012b03,
		32'h02010113,
		32'h00008067,
		32'h00002537,
		32'h92050513,
		32'hf18ff0ef,
		32'h00400793,
		32'hfc1ff06f,
		32'hfff00513,
		32'hfc1ff06f,
		32'hfe010113,
		32'h00812c23,
		32'h00912a23,
		32'h01212823,
		32'h01312623,
		32'h01412423,
		32'h01512223,
		32'h00112e23,
		32'h00050993,
		32'h00058a13,
		32'h00060413,
		32'h00068493,
		32'h00070913,
		32'hfff00a93,
		32'h9c9ff0ef,
		32'h05551663,
		32'h00048693,
		32'h00040613,
		32'h000a0593,
		32'h00098513,
		32'hdd1ff0ef,
		32'h03551a63,
		32'h00040513,
		32'h01812403,
		32'h01c12083,
		32'h00c12983,
		32'h00812a03,
		32'h00412a83,
		32'h00090613,
		32'h00048593,
		32'h01012903,
		32'h01412483,
		32'h02010113,
		32'hbedff06f,
		32'h01c12083,
		32'h01812403,
		32'h01412483,
		32'h01012903,
		32'h00c12983,
		32'h00812a03,
		32'h00412a83,
		32'h02010113,
		32'h00008067,
		32'he5010113,
		32'h1a812423,
		32'h1a912223,
		32'h19312e23,
		32'h19412c23,
		32'h1a112623,
		32'h1b212023,
		32'h19512a23,
		32'h00050493,
		32'h00058a13,
		32'h00060993,
		32'h00068413,
		32'h80001737,
		32'h80c72783,
		32'hfe079ee3,
		32'h19000613,
		32'h00000593,
		32'h00010513,
		32'hf08ff0ef,
		32'h8c1647b7,
		32'h54978793,
		32'h00f12023,
		32'h25ac97b7,
		32'hc1678793,
		32'h00f12223,
		32'h454927b7,
		32'h50178793,
		32'h00f12423,
		32'h000047b7,
		32'h50078793,
		32'h00f12623,
		32'h400047b7,
		32'h00678793,
		32'h00f12a23,
		32'h0000d7b7,
		32'hac578793,
		32'h00f12c23,
		32'h0f8107b7,
		32'h00f12e23,
		32'h000067b7,
		32'h02f12623,
		32'hfaf007b7,
		32'h02f12823,
		32'h20400793,
		32'h02f12a23,
		32'h05b407b7,
		32'h02f12c23,
		32'h01c4d783,
		32'h0104a703,
		32'h00c00593,
		32'h00f11e23,
		32'h01e4d783,
		32'h00c10513,
		32'h05a40913,
		32'h02f11123,
		32'h000027b7,
		32'h70778793,
		32'h00f707b3,
		32'h00170713,
		32'h00f11823,
		32'h00e4a823,
		32'h02c40793,
		32'h00f11923,
		32'hc3dff0ef,
		32'h00050a93,
		32'h14040a63,
		32'h0009c783,
		32'h0019c703,
		32'h00010693,
		32'h00879793,
		32'h00e7e7b3,
		32'h02f11c23,
		32'h00298713,
		32'h413707b3,
		32'h00468693,
		32'h0e87cc63,
		32'h00180737,
		32'h01041793,
		32'h00670713,
		32'h00e787b3,
		32'h40145413,
		32'h00f12a23,
		32'h01440593,
		32'h0264d783,
		32'h01410513,
		32'h02f11023,
		32'h01a4d783,
		32'h02f11323,
		32'h0084d783,
		32'h02f11223,
		32'h00a4d783,
		32'h02f11523,
		32'h00c4d783,
		32'h02f11423,
		32'h00e4d783,
		32'h02f11723,
		32'h02c15783,
		32'h00fa6a33,
		32'h03411623,
		32'hbadff0ef,
		32'h000047b7,
		32'h00f11b23,
		32'h04000793,
		32'h00f10aa3,
		32'h000017b7,
		32'h80078793,
		32'h80001737,
		32'h800016b7,
		32'h00f11723,
		32'h02a11823,
		32'h01511d23,
		32'h00010793,
		32'h82070713,
		32'h9b068613,
		32'h0007a583,
		32'h00470713,
		32'h00478793,
		32'hfeb72e23,
		32'hfec718e3,
		32'h8126a023,
		32'h8006a223,
		32'h8006a423,
		32'h00300793,
		32'h00002537,
		32'h84850513,
		32'h80f6a623,
		32'hc60ff0ef,
		32'h1ac12083,
		32'h1a812403,
		32'h1a412483,
		32'h1a012903,
		32'h19c12983,
		32'h19812a03,
		32'h19412a83,
		32'h00000513,
		32'h1b010113,
		32'h00008067,
		32'h00074783,
		32'h00174603,
		32'h00470713,
		32'h01879793,
		32'h01061613,
		32'h00c7e7b3,
		32'hfff74603,
		32'h00c7e7b3,
		32'hffe74603,
		32'h00861613,
		32'h00c7e7b3,
		32'h02f6ac23,
		32'hed1ff06f,
		32'h001807b7,
		32'h00678793,
		32'h00f12a23,
		32'h01400593,
		32'hee5ff06f,
		32'hfc010113,
		32'h02912a23,
		32'h03412423,
		32'h800004b7,
		32'h10000a37,
		32'h02812c23,
		32'h03212823,
		32'h03312623,
		32'h03512223,
		32'h03612023,
		32'h01712e23,
		32'h01812c23,
		32'h01912a23,
		32'h01a12823,
		32'h01b12623,
		32'h02112e23,
		32'h00050413,
		32'h00058993,
		32'h00060d93,
		32'h00c48913,
		32'h02650a93,
		32'h02850b13,
		32'h02050b93,
		32'h01c50c13,
		32'h01450c93,
		32'h017a0d13,
		32'h00100793,
		32'h00092703,
		32'hfef71ee3,
		32'h000a8713,
		32'h000b0693,
		32'h000b8613,
		32'h000c0593,
		32'h000c8513,
		32'hc61ff0ef,
		32'h01a57733,
		32'h0149e7b3,
		32'h12f71263,
		32'h04c4d703,
		32'h0324d483,
		32'h00a75793,
		32'h40f484b3,
		32'hfec48493,
		32'h0a049663,
		32'h00357793,
		32'h0e079e63,
		32'h80000737,
		32'h04475783,
		32'h04a75603,
		32'h01079793,
		32'h00c787b3,
		32'h009787b3,
		32'h0107d613,
		32'h00c41623,
		32'h00f41723,
		32'h04875783,
		32'h00f41423,
		32'h04e75783,
		32'h00f41523,
		32'h100007b7,
		32'h00278793,
		32'h00f51c63,
		32'h04075783,
		32'h00f41d23,
		32'h567817b7,
		32'h23478793,
		32'h00f42423,
		32'h80000537,
		32'h00c50513,
		32'h8c9ff0ef,
		32'h03c12083,
		32'h03812403,
		32'h03012903,
		32'h02c12983,
		32'h02812a03,
		32'h02412a83,
		32'h02012b03,
		32'h01c12b83,
		32'h01812c03,
		32'h01412c83,
		32'h01012d03,
		32'h00c12d83,
		32'h00048513,
		32'h03412483,
		32'h04010113,
		32'h00008067,
		32'h00c75793,
		32'h00e78793,
		32'h00279793,
		32'h012787b3,
		32'hffd7c703,
		32'h00ed8023,
		32'hffc7c703,
		32'h00ed80a3,
		32'h002d8713,
		32'h41b706b3,
		32'hf296d8e3,
		32'h0037c683,
		32'h00470713,
		32'h00478793,
		32'hfed70e23,
		32'hffe7c683,
		32'hfed70ea3,
		32'hffd7c683,
		32'hfed70f23,
		32'hffc7c683,
		32'hfed70fa3,
		32'hfd1ff06f,
		32'h00100493,
		32'hf05ff06f,
		32'h00090513,
		32'h821ff0ef,
		32'hea9ff06f,
		32'h6cbe57b7,
		32'h60278793,
		32'h00f52423,
		32'h454997b7,
		32'hc1678793,
		32'h02f52023,
		32'haf5127b7,
		32'h50178793,
		32'h02f52223,
		32'h0f81d7b7,
		32'hac578793,
		32'h00b52023,
		32'h00052223,
		32'h00052623,
		32'h00052823,
		32'h02f52423,
		32'h00008067,
		32'h0065d783,
		32'hfe010113,
		32'h00112e23,
		32'h00812c23,
		32'h00f51d23,
		32'h0085d783,
		32'h00000693,
		32'h00c10613,
		32'h00f51e23,
		32'h00a5d783,
		32'h00200593,
		32'h00050413,
		32'h00f51f23,
		32'h454997b7,
		32'hc1678793,
		32'h00f52a23,
		32'h000027b7,
		32'h5ac78793,
		32'h00f51c23,
		32'hb41ff0ef,
		32'h00c10613,
		32'h01200593,
		32'h00040513,
		32'hd9dff0ef,
		32'h00c10613,
		32'h00040513,
		32'h00000693,
		32'h01000593,
		32'hb1dff0ef,
		32'h01c12083,
		32'h01812403,
		32'h02010113,
		32'h00008067,
		32'h0125d783,
		32'h02f51323,
		32'h0145d783,
		32'h02f51423,
		32'h0165d783,
		32'h02f51523,
		32'h00008067,
		32'hfe010113,
		32'h00812c23,
		32'h00c10613,
		32'h00058413,
		32'h00200593,
		32'h00112e23,
		32'h00912a23,
		32'h00050493,
		32'hd39ff0ef,
		32'h00c10613,
		32'h00000693,
		32'h01200593,
		32'h00048513,
		32'hab9ff0ef,
		32'h00040513,
		32'h924ff0ef,
		32'h01c12083,
		32'h01812403,
		32'h01412483,
		32'h02010113,
		32'h00008067,
		32'hfe010113,
		32'h00812c23,
		32'h00c10613,
		32'h00058413,
		32'h01000593,
		32'h00912a23,
		32'h00112e23,
		32'h00050493,
		32'hce5ff0ef,
		32'h0004a783,
		32'h00f42023,
		32'h0044a783,
		32'h00f42223,
		32'h0084d783,
		32'h00f41423,
		32'h00a4d783,
		32'h00f41523,
		32'h00c4d783,
		32'h00f41623,
		32'h00e4d783,
		32'h00f41723,
		32'h0104a783,
		32'h00f42823,
		32'h0144d783,
		32'h00f41a23,
		32'h0164d783,
		32'h00f41b23,
		32'h0184d783,
		32'h00f41c23,
		32'h01a4d783,
		32'h00f41d23,
		32'h01c4d783,
		32'h00f41e23,
		32'h01e4d783,
		32'h00f41f23,
		32'h0204d783,
		32'h02f41023,
		32'h0224d783,
		32'h02f41123,
		32'h0244d783,
		32'h02f41223,
		32'h0264d783,
		32'h01c12083,
		32'h02f41323,
		32'h0284d783,
		32'h02f41423,
		32'h02a4d783,
		32'h01412483,
		32'h02f41523,
		32'h01812403,
		32'h02010113,
		32'h00008067,
		32'h00052783,
		32'hff010113,
		32'h00112623,
		32'h00812423,
		32'h00912223,
		32'h04079263,
		32'h00058493,
		32'h00060693,
		32'h00058613,
		32'h01000593,
		32'h00050413,
		32'h99dff0ef,
		32'h00048613,
		32'h01000593,
		32'h00040513,
		32'hbf9ff0ef,
		32'h00c12083,
		32'h00812403,
		32'h00412483,
		32'h00000513,
		32'h01010113,
		32'h00008067,
		32'h0f0000ef,
		32'hfe5ff06f,
		32'h00052783,
		32'hfc010113,
		32'h02912a23,
		32'h02112e23,
		32'h02812c23,
		32'h03212823,
		32'h03312623,
		32'h00060493,
		32'h04079c63,
		32'h00058613,
		32'h00058993,
		32'h01000593,
		32'h00050913,
		32'hba1ff0ef,
		32'h00050413,
		32'h00000693,
		32'h00098613,
		32'h01000593,
		32'h00090513,
		32'h91dff0ef,
		32'h00040513,
		32'h0084d463,
		32'h00048513,
		32'h03c12083,
		32'h03812403,
		32'h03412483,
		32'h03012903,
		32'h02c12983,
		32'h04010113,
		32'h00008067,
		32'h00810613,
		32'h288000ef,
		32'h00050413,
		32'hfcdff06f,
		32'h00052783,
		32'h04079c63,
		32'hfe010113,
		32'h00000693,
		32'h00c10613,
		32'h01100593,
		32'h00112e23,
		32'h00812c23,
		32'h00050413,
		32'h8bdff0ef,
		32'h00c10613,
		32'h01100593,
		32'h00040513,
		32'hb19ff0ef,
		32'h00c10613,
		32'h00040513,
		32'h00000693,
		32'h01000593,
		32'h899ff0ef,
		32'h01c12083,
		32'h01812403,
		32'h02010113,
		32'h00008067,
		32'h00008067,
		32'he5010113,
		32'h1a812423,
		32'h1a912223,
		32'h19412c23,
		32'h1a112623,
		32'h1b212023,
		32'h19312e23,
		32'h19512a23,
		32'h19612823,
		32'h00050493,
		32'h00058a13,
		32'h00060413,
		32'h80001737,
		32'h80c72783,
		32'hfe079ee3,
		32'h19000613,
		32'h00000593,
		32'h00010513,
		32'hf89fe0ef,
		32'h8c1647b7,
		32'h54978793,
		32'h00f12023,
		32'h25ac97b7,
		32'hc1678793,
		32'h00f12223,
		32'h454927b7,
		32'h50178793,
		32'h00f12423,
		32'h000047b7,
		32'h50078793,
		32'h00f12623,
		32'h400047b7,
		32'h01178793,
		32'h00f12a23,
		32'h0000d7b7,
		32'hac578793,
		32'h00f12c23,
		32'h0f8107b7,
		32'h00f12e23,
		32'h01c4d783,
		32'h0104a703,
		32'h01041a93,
		32'h00f11e23,
		32'h01e4d783,
		32'h010ada93,
		32'h00c00593,
		32'h02f11123,
		32'h000027b7,
		32'h70778793,
		32'h00f707b3,
		32'h00170713,
		32'h00f11823,
		32'h00e4a823,
		32'h01ca8793,
		32'h00c10513,
		32'h00f11923,
		32'hcd8ff0ef,
		32'h000a4783,
		32'h001a4703,
		32'h00010913,
		32'h00879793,
		32'h00e7e7b3,
		32'h04a40993,
		32'h00050b13,
		32'h02f11423,
		32'h002a0713,
		32'h00090693,
		32'h414707b3,
		32'h00468693,
		32'h0c87ca63,
		32'h00080737,
		32'h01170713,
		32'h01041793,
		32'h00e787b3,
		32'h00f12a23,
		32'h0264d783,
		32'h40145593,
		32'h008a8a93,
		32'h02f11023,
		32'h01a4d783,
		32'h01058593,
		32'h01410513,
		32'h02f11323,
		32'h03511223,
		32'hc68ff0ef,
		32'h000047b7,
		32'h00f11b23,
		32'h04000793,
		32'h00f10aa3,
		32'h000017b7,
		32'h80078793,
		32'h00f11723,
		32'h80001737,
		32'h800017b7,
		32'h02a11523,
		32'h01611d23,
		32'h82078793,
		32'h9b070693,
		32'h00092603,
		32'h00478793,
		32'h00490913,
		32'hfec7ae23,
		32'hfed798e3,
		32'h81372023,
		32'h80072223,
		32'h80072423,
		32'h00300793,
		32'h00002537,
		32'h84850513,
		32'h80f72623,
		32'hd21fe0ef,
		32'h1ac12083,
		32'h1a812403,
		32'h1a412483,
		32'h1a012903,
		32'h19c12983,
		32'h19812a03,
		32'h19412a83,
		32'h19012b03,
		32'h00000513,
		32'h1b010113,
		32'h00008067,
		32'h00074783,
		32'h00174603,
		32'h00470713,
		32'h01879793,
		32'h01061613,
		32'h00c7e7b3,
		32'hfff74603,
		32'h00c7e7b3,
		32'hffe74603,
		32'h00861613,
		32'h00c7e7b3,
		32'h02f6a423,
		32'hef5ff06f,
		32'hfd010113,
		32'h01312e23,
		32'h800009b7,
		32'h02812423,
		32'h02912223,
		32'h03212023,
		32'h01412c23,
		32'h01512a23,
		32'h01612823,
		32'h01712623,
		32'h01812423,
		32'h01912223,
		32'h01a12023,
		32'h02112623,
		32'h00058413,
		32'h00060913,
		32'h00100a93,
		32'h00c98a13,
		32'h02650b13,
		32'h02850b93,
		32'h02050c13,
		32'h01c50c93,
		32'h01450493,
		32'h20000d37,
		32'h000a2783,
		32'hff579ee3,
		32'h000b0713,
		32'h000b8693,
		32'h000c0613,
		32'h000c8593,
		32'h00048513,
		32'hd3cff0ef,
		32'h0ba51e63,
		32'h0409d703,
		32'h00240593,
		32'h800006b7,
		32'h00e91323,
		32'h0389d703,
		32'h00e91423,
		32'h03e9d783,
		32'h00f91523,
		32'h0499c783,
		32'h0449d483,
		32'h00f40023,
		32'h0489c783,
		32'hff848493,
		32'h00f400a3,
		32'h00200793,
		32'h0497c663,
		32'h80000537,
		32'h00c50513,
		32'h9e0ff0ef,
		32'h02c12083,
		32'h02812403,
		32'h02012903,
		32'h01c12983,
		32'h01812a03,
		32'h01412a83,
		32'h01012b03,
		32'h00c12b83,
		32'h00812c03,
		32'h00412c83,
		32'h00012d03,
		32'h00048513,
		32'h02412483,
		32'h03010113,
		32'h00008067,
		32'h00f68733,
		32'h04d74603,
		32'h00478793,
		32'h00458593,
		32'hfec58e23,
		32'h04c74603,
		32'hfec58ea3,
		32'h04b74603,
		32'hfec58f23,
		32'h04a74703,
		32'hfee58fa3,
		32'hf89ff06f,
		32'h000a0513,
		32'h96cff0ef,
		32'hf1dff06f,
		32'h0065d783,
		32'h00f51d23,
		32'h0085d783,
		32'h00f51e23,
		32'h00a5d783,
		32'h00f51f23,
		32'h000027b7,
		32'h5ac78793,
		32'h00f51a23,
		32'h00100513,
		32'h00008067,
		32'hfe010113,
		32'h00912a23,
		32'h00058493,
		32'h00068593,
		32'h00812c23,
		32'h00c12623,
		32'h00112e23,
		32'h00050413,
		32'hfb5ff0ef,
		32'h00c12603,
		32'h00100793,
		32'hfff00513,
		32'h00c7da63,
		32'h00048593,
		32'h00040513,
		32'hc35ff0ef,
		32'h00000513,
		32'h01c12083,
		32'h01812403,
		32'h01412483,
		32'h02010113,
		32'h00008067,
		32'hff010113,
		32'h00812423,
		32'h00060413,
		32'h00068613,
		32'h00112623,
		32'he21ff0ef,
		32'h00a45463,
		32'h00040513,
		32'h00c12083,
		32'h00812403,
		32'h01010113,
		32'h00008067,
		32'h06054063,
		32'h0605c663,
		32'h00058613,
		32'h00050593,
		32'hfff00513,
		32'h02060c63,
		32'h00100693,
		32'h00b67a63,
		32'h00c05863,
		32'h00161613,
		32'h00169693,
		32'hfeb66ae3,
		32'h00000513,
		32'h00c5e663,
		32'h40c585b3,
		32'h00d56533,
		32'h0016d693,
		32'h00165613,
		32'hfe0696e3,
		32'h00008067,
		32'h00008293,
		32'hfb5ff0ef,
		32'h00058513,
		32'h00028067,
		32'h40a00533,
		32'h0005d863,
		32'h40b005b3,
		32'hf9dff06f,
		32'h40b005b3,
		32'h00008293,
		32'hf91ff0ef,
		32'h40a00533,
		32'h00028067,
		32'h00008293,
		32'h0005ca63,
		32'h00054c63,
		32'hf79ff0ef,
		32'h00058513,
		32'h00028067,
		32'h40b005b3,
		32'hfe0558e3,
		32'h40a00533,
		32'hf61ff0ef,
		32'h40b00533,
		32'h00028067,
		32'h00001941,
		32'h73697200,
		32'h01007663,
		32'h0000000f,
		32'h33767205,
		32'h70326932,
		32'h00000030,
		32'h73654d0a,
		32'h65676173,
		32'h6f726620,
		32'h6573206d,
		32'h72657672,
		32'h0000203a,
		32'h202c6948,
		32'h206d2749,
		32'h75546f41,
		32'h216e616d,
		32'h0000000a,
		32'h00000000,
		32'h00000000,
		32'h00000000,
		32'h00000000,
		32'h00000000,
		32'h3a434347,
		32'h4e472820,
		32'h39202955,
		32'h302e322e,
		32'h001b4100,
		32'h69720000,
		32'h00766373,
		32'h00001101,
		32'h05100400,
		32'h32337672,
		32'h30703269,
		32'h00000000,
		32'h33323130,
		32'h37363534,
		32'h42413938,
		32'h46454443,
		32'h00000000,
		32'h696e6946,
		32'h0a216873,
		32'h001b4100,
		32'h69720000,
		32'h00766373,
		32'h00001101,
		32'h05100400,
		32'h32337672,
		32'h30703269,
		32'h00000000,
		32'h646e6553,
		32'h70726120,
		32'h00000a21,
		32'h76636552,
		32'h50524120,
		32'h7165522d,
		32'h6e61202c,
		32'h65732064,
		32'h4120646e,
		32'h522d5052,
		32'h21707365,
		32'h0000000a,
		32'h76636552,
		32'h50524120,
		32'h7365522d,
		32'h000a2170,
		32'h646e6573,
		32'h6d636920,
		32'h65722070,
		32'h75732071,
		32'h73656363,
		32'h6c756673,
		32'h000a796c,
		32'h75746552,
		32'h69206e72,
		32'h20706d63,
		32'h70736572,
		32'h63757320,
		32'h73736563,
		32'h6c6c7566,
		32'h000a2179,
		32'h63736964,
		32'h20647261,
		32'h6b636170,
		32'h000a7465,
		32'h3d3d3d0a,
		32'h3d3d3d3d,
		32'h3d3d3d3d,
		32'h3d3d3d3d,
		32'h00000a3d,
		32'h646e6573,
		32'h0000000a,
		32'h76636572,
		32'h6d636920,
		32'h65722070,
		32'h000a2171,
		32'h76636572,
		32'h6d636920,
		32'h65722070,
		32'h0a217073,
		32'h00000000,
		32'hffffffff,
		32'hffff0000,
		32'h00000000,
		32'h08060001,
		32'h08000604,
		32'h00010000,
		32'h00000000,
		32'hcac50f81,
		32'h00000000,
		32'h00000000,
		32'h00000000,
		32'h00000000,
		32'h00000000,
		32'h00000000,
		32'h00000000,
		32'h00000000,
		32'h0000004a,
		32'h00000000,
		32'h00000000,
		32'h00000003,
		32'h00000000,
		32'h00000000,
		32'h00000000,
		32'h08004500,
		32'h00542baf,
		32'h40004001,
		32'h5a6c0000,
		32'h00000000,
		32'h00000800,
		32'hf961500b,
		32'h0001bdd4,
		32'h365e0000,
		32'h0000f28b,
		32'h09000000,
		32'h00001011,
		32'h12131415,
		32'h16171819,
		32'h1a1b1c1d,
		32'h1e1f2021,
		32'h22232425,
		32'h26272829,
		32'h2a2b2c2d,
		32'h2e2f3031,
		32'h32333435,
		32'h36370000,
		32'h00000000,
		32'h00000000,
		32'h00000000,
		32'h00000082,
		32'h00000000,
		32'h00000000,
		32'h00000003,
		32'h00001b41,
		32'h73697200,
		32'h01007663,
		32'h00000011,
		32'h72051004,
		32'h69323376,
		32'h00307032,
		32'h00001b41,
		32'h73697200,
		32'h01007663,
		32'h00000011,
		32'h72051004,
		32'h69323376,
		32'h00307032,
		32'h00001b41,
		32'h73697200,
		32'h01007663,
		32'h00000011,
		32'h72051004,
		32'h69323376,
		32'h00307032,
		32'h00001941,
		32'h73697200,
		32'h01007663,
		32'h0000000f,
		32'h33767205,
		32'h70326932,
		32'h00000030,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0,
		32'h0
    };

	// reg 	[31:0] 	memory [0:64*1024/4-1];
	
	reg 	[13:0] 	addr_q;
    wire 	[31:0]	memory_data;
    reg 	[31:0]	addr_conf;

    reg 	[3:0]	count,pkt_count;

     always @* begin
    	addr_q <= 13'h7ff - addr_conf[10:0];
    end
	assign memory_data = memory[addr_q];

	reg [4:0]	state_mem;
	parameter 	IDLE_S 		= 5'd0,
				FAKE_DATA_S	= 5'd1,
				CONF_TCM_S	= 5'd2,
				CONF_TCM_1_S= 5'd3,
				CONF_TCM_2_S= 5'd4,
				CONF_SEL_1_S= 5'd5,
				CONF_SEL_2_S= 5'd6,
				READY_S		= 5'd7,
				READ_1_S	= 5'd8,
				READ_2_S	= 5'd9,
				READ_3_S	= 5'd10,
				READ_4_S	= 5'd11,
				READ_5_S	= 5'd12,
				READ_6_S	= 5'd13,
				WRITE_END_S	= 5'd14,
				WAIT_10_CLK_S= 5'd15,
				TEST_L2SW_S	= 5'd16;

	always @(posedge clk or negedge resetn) begin
		if (!resetn) begin
			// reset
//			addr_q 		<= 14'h400;
			state_mem 	<= IDLE_S;

			data_in_valid	<= 1'b0;
			data_in 		<= 134'b0;
			count			<= 4'b0;
			pkt_count		<= 4'b0;
			addr_conf		<= 32'b0;
		end
		else begin
			case(state_mem)
				IDLE_S: begin
					data_in_valid 	<= 1'b1;
					data_in 		<= {2'b01,4'b0,128'b0};
					state_mem 		<= FAKE_DATA_S;
					count 			<= 4'b0;
				end
				FAKE_DATA_S: begin
					count <= count + 4'd1;
					case(count)
						4'd0: data_in <= {2'b11, 4'b0, 128'd0};
						4'd1: data_in <= {2'b11, 4'b0, 96'b0,16'h9001,16'b0};
						4'd2: data_in <= {2'b11, 4'b0, 112'd1,16'b0};
						4'd3: data_in <= {2'b11, 4'b0, 112'd2,16'b0};
						4'd4: data_in <= {2'b11, 4'b0, 112'd3,16'b0};
						4'd5: data_in <= {2'b10, 4'b0, 112'd4,16'b0};
						default: begin
						end
					endcase
					if(count == 4'd5)
						state_mem <= CONF_TCM_S;
				end
				CONF_TCM_S: begin
					data_in_valid 	<= 1'b1;
					data_in 		<= {2'b01,4'b0,128'b0};
					state_mem 		<= CONF_TCM_1_S;
					count 			<= 4'b0;
				end
				CONF_TCM_1_S: begin
					count <= count + 4'd1;
					case(count)
						4'd0: data_in <= {2'b11, 4'b0, 128'd0};
						4'd1: data_in <= {2'b11, 4'b0, 96'b0,16'h9003,16'b0};
						default: begin
						end
					endcase
					if(count == 4'd1)
						state_mem <= CONF_TCM_2_S;
					//addr_q <= 14'h3ff;
					addr_conf <= 32'b0;
				end
				CONF_TCM_2_S: begin
					addr_conf 	<= addr_conf + 32'd1;
					//addr_q 		<= addr_q - 14'd1;
					data_in[131:0] <= {4'b0, 48'd0, memory_data, addr_conf,16'b0};
					if(addr_conf == 32'd2000) begin
						state_mem <= READ_1_S;
						data_in[133:132] <= {2'b10};
					end
					else begin
						state_mem <= CONF_TCM_2_S;
						data_in[133:132] <= {2'b11};
					end
				end
				CONF_SEL_1_S: begin
					data_in_valid 	<= 1'b1;
					data_in 		<= {2'b01,4'b0,128'b0};
					state_mem 		<= CONF_SEL_2_S;
					count 			<= 4'b0;
				end
				CONF_SEL_2_S: begin
					count <= count + 4'd1;
					case(count)
						4'd0: data_in <= {2'b11, 4'b0, 128'd0};
						4'd1: data_in <= {2'b11, 4'b0, 96'b0,16'h9001,16'b0};
						4'd2: data_in <= {2'b11, 4'b0, 128'd0};
						4'd3: data_in <= {2'b11, 4'b0, 128'd1};
						4'd4: data_in <= {2'b11, 4'b0, 128'd2};
						4'd5: data_in <= {2'b10, 4'b0, 128'd3};
						default: begin
						end
					endcase
					if(count == 4'd5) begin
						count		<= 4'd0;
						// state_mem 	<= WAIT_10_CLK_S;
						state_mem 	<= READY_S;
					end
				end
				READ_1_S: begin
					data_in_valid 	<= 1'b1;
					data_in 		<= {2'b01,4'b0,128'b0};
					state_mem 		<= READ_2_S;
					count 			<= 4'b0;
				end
				READ_2_S: begin
					count <= count + 4'd1;
					case(count)
						4'd0: data_in <= {2'b11, 4'b0, 128'd0};
						4'd1: data_in <= {2'b11, 4'b0, 96'b0,16'h9002,16'b0};
						4'd2: data_in <= {2'b11, 4'b0, 128'd1};
						4'd3: data_in <= {2'b11, 4'b0, 128'd2};
						4'd4: data_in <= {2'b11, 4'b0, 128'd3};
						4'd5: data_in <= {2'b10, 4'b0, 128'd4};
						default: begin
						end
					endcase
					if(count == 4'd5)
						state_mem <= READ_3_S;
				end
				READ_3_S: begin
					data_in_valid 	<= 1'b1;
					data_in 		<= {2'b01,4'b0,128'b0};
					state_mem 		<= READ_4_S;
					count 			<= 4'b0;
				end
				READ_4_S: begin
					count <= count + 4'd1;
					case(count)
						4'd0: data_in <= {2'b11, 4'b0, 128'd0};
						4'd1: data_in <= {2'b11, 4'b0, 96'b0,16'h9004,16'b0};
						4'd2: data_in <= {2'b11, 4'b0, 112'd128,16'b0};
						4'd3: data_in <= {2'b11, 4'b0, 128'd2};
						4'd4: data_in <= {2'b11, 4'b0, 128'd3};
						4'd5: data_in <= {2'b10, 4'b0, 128'd4};
						default: begin
						end
					endcase
					if(count == 4'd5)
						state_mem <= READ_5_S;
				end
				READ_5_S: begin
					data_in_valid 	<= 1'b1;
					data_in 		<= {2'b01,4'b0,128'b0};
					state_mem 		<= READ_6_S;
					count 			<= 4'b0;
				end
				READ_6_S: begin
					count <= count + 4'd1;
					case(count)
						4'd0: data_in <= {2'b11, 4'b0, 128'd0};
						4'd1: data_in <= {2'b11, 4'b0, 96'b0,16'h9004,16'b0};
						4'd2: data_in <= {2'b11, 4'b0, 112'd129,16'b0};
						4'd3: data_in <= {2'b11, 4'b0, 128'd2};
						4'd4: data_in <= {2'b11, 4'b0, 128'd3};
						4'd5: data_in <= {2'b10, 4'b0, 128'd4};
						default: begin
						end
					endcase
					if(count == 4'd5)
						state_mem <= CONF_SEL_1_S;
				end
				WAIT_10_CLK_S: begin
					data_in_valid		<= 1'b0;
					count 				<= count + 4'd1;
					if(count == 4'd10) begin
						count 			<= 4'd0;
						data_in_valid 	<= 1'b1;
						data_in 		<= {2'b01,4'b0,128'b0};
						state_mem		<= TEST_L2SW_S;
					end
					else 
						state_mem		<= WAIT_10_CLK_S;
				end
				TEST_L2SW_S: begin
					count <= count + 4'd1;
					case(count)
						4'd0: data_in <= {2'b11, 4'b0, 128'd0};
						4'd1: data_in <= {2'b11, 4'b0, 48'hffff_ffff_ffff, 48'b0,16'h0800,16'b0};
						4'd2: data_in <= {2'b11, 4'b0, 64'd6,64'd0};
						4'd3: data_in <= {2'b11, 4'b0, 128'd1};
						4'd4: data_in <= {2'b11, 4'b0, 128'd2};
						4'd5: data_in <= {2'b10, 4'b0, 128'd3};
						default: begin
						end
					endcase
					if(count == 4'd5) begin
						count			<= 4'd0;
						if(pkt_count == 4'd4)
							state_mem	<= READY_S;
						else begin
							state_mem 	<= WAIT_10_CLK_S;
							pkt_count	<= 4'd1 + pkt_count;
						end
					end
				end
				READY_S: begin
					data_in_valid <= 1'b0;
					state_mem <= READY_S;
				end
				default: begin
					state_mem <= IDLE_S;
				end
			endcase
		end
	end


endmodule
