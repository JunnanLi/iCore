/*
 *  iCore_hardware -- Hardware for TuMan RISC-V (RV32I) Processor Core.
 *
 *  Copyright (C) 2019-2020 Junnan Li <lijunnan@nudt.edu.cn>.
 *  Copyright and related rights are licensed under the MIT license.
 *
 *	Data: 2020.01.01
 *	Description: This module is used to connect TuMan_top and configuration.
 */

/**	Please toggle following comment (i.e., `define FPGA_ALTERA) if you 
 **	 use an Alater (Intel) FPGA
 **/
// `define FPGA_ALTERA

module um_for_cpu(
	input				clk,
	input				rst_n,
    
	// FAST packets from CPU (ARM A8) or Physical ports, the format is according to fast 
	//	 project (www.http://www.fastswitch.org/)
	input				data_in_valid,
	input		[133:0] data_in,	// 2'b01 is head, 2'b00 is body, and 2'b10 is tail;
	
	output reg			data_out_valid,
	output reg	[133:0] data_out,
	output wire			mem_wren,
	output wire			mem_rden,
	output wire	[31:0]	mem_addr,
	output wire	[31:0]	mem_wdata,
	input		[31:0]	mem_rdata,
	output wire			cpu_ready
);

	/**	TODO:*/

	wire 		conf_rden_itcm, conf_wren_itcm, conf_rden_dtcm, conf_wren_dtcm;
	wire [31:0]	conf_addr_itcm, conf_wdata_itcm, conf_rdata_itcm;
	wire [31:0]	conf_addr_dtcm, conf_wdata_dtcm, conf_rdata_dtcm;
	wire 		conf_sel_dtcm;
	wire 		print_valid;
	wire [7:0]	print_value;
	wire		data_valid_confMem;
	wire [133:0]data_confMem;
	// fifo interface
	reg			rdreq_pkt;
	wire [133:0]q_pkt;
	reg	 [7:0]	count_pkt;	// number of packet in the fifo;
	
	assign cpu_ready= ~conf_sel_dtcm;

	TuMan32_top tm(
		.clk(clk),
		.resetn(rst_n),

		.conf_rden_itcm(conf_rden_itcm),
		.conf_wren_itcm(conf_wren_itcm),
		.conf_addr_itcm(conf_addr_itcm),
		.conf_wdata_itcm(conf_wdata_itcm),
		.conf_rdata_itcm(conf_rdata_itcm),

		.conf_sel_dtcm(conf_sel_dtcm),
		.conf_rden_dtcm(conf_rden_dtcm),
		.conf_wren_dtcm(conf_wren_dtcm),
		.conf_addr_dtcm(conf_addr_dtcm),
		.conf_wdata_dtcm(conf_wdata_dtcm),
		.conf_rdata_dtcm(conf_rdata_dtcm),

		.print_valid(print_valid),
		.print_value(print_value),

		.mem_wren_toPipe(mem_wren),
		.mem_rden_toPipe(mem_rden),
		.mem_addr_toPipe(mem_addr),
		.mem_wdata_toPipe(mem_wdata),
		.mem_rdata_fromPipe(mem_rdata)
	);

	conf_mem confMem(
		.clk(clk),
		.resetn(rst_n),

		.data_in_valid(data_in_valid),
		.data_in(data_in),
		.data_out_valid(data_valid_confMem),
		.data_out(data_confMem),

		.conf_rden_itcm(conf_rden_itcm),
		.conf_wren_itcm(conf_wren_itcm),
		.conf_addr_itcm(conf_addr_itcm),
		.conf_wdata_itcm(conf_wdata_itcm),
		.conf_rdata_itcm(conf_rdata_itcm),

		.conf_sel_dtcm(conf_sel_dtcm),
		.conf_rden_dtcm(conf_rden_dtcm),
		.conf_wren_dtcm(conf_wren_dtcm),
		.conf_addr_dtcm(conf_addr_dtcm),
		.conf_wdata_dtcm(conf_wdata_dtcm),
		.conf_rdata_dtcm(conf_rdata_dtcm),

		.print_valid(print_valid),
		.print_value(print_value)
	);


	/**	fifo used to store packet generated by cpu*/
`ifdef FPGA_ALTERA
	fifo pkt_buffer(
		.aclr(!rst_n),
		.clock(clk),
		.data(data_confMem),
		.rdreq(rdreq_pkt),
		.wrreq(data_valid_confMem),
		.empty(),
		.full(),
		.q(q_pkt),
		.usedw()
	);
	defparam
		pkt_buffer.width = 134,
		pkt_buffer.depth = 9,
		pkt_buffer.words = 256;
`else
	fifo_134_512 pkt_buffer(
		.clk(clk),
		.srst(!rst_n),
		.din(data_confMem),
		.wr_en(data_valid_confMem),
		.rd_en(rdreq_pkt),
		.dout(q_pkt),
		.full(),
		.empty()
	);
`endif

	/** output packet */
	reg			state_out;
	parameter	IDLE_S		= 1'b0,
				READ_FIFO_S	= 1'b1;
	always @(posedge clk or negedge rst_n) begin
		if (!rst_n) begin
			// reset
			count_pkt		<= 8'b0;
			// output packet;
			state_out		<= IDLE_S;
			data_out_valid	<= 1'b0;
			data_out		<= 134'b0;
			rdreq_pkt		<= 1'b0;
		end
		else begin
			if((data_confMem[133:132] == 2'b10 && data_valid_confMem == 1'b1) &&
				(data_out[133:132] == 2'b01 && data_out_valid == 1'b1))
					count_pkt	<= count_pkt;
			else if(data_confMem[133:132] == 2'b10 && data_valid_confMem == 1'b1)
				count_pkt		<= count_pkt + 8'd1;
			else if(data_out[133:132] == 2'b01 && data_out_valid == 1'b1)
				count_pkt		<= count_pkt - 8'd1;
			else
				count_pkt		<= count_pkt;

			(* full_case *)
			case(state_out)
				IDLE_S: begin
					data_out_valid	<= 1'b0;
					if(count_pkt != 0) begin
						rdreq_pkt	<= 1'b1;
						state_out	<= READ_FIFO_S;
					end
					else begin
						rdreq_pkt	<= 1'b0;
						state_out	<= IDLE_S;
					end
				end
				READ_FIFO_S: begin
					data_out_valid	<= 1'b1;
					data_out		<= q_pkt;
					if(q_pkt[133:132] == 2'b10) begin
						rdreq_pkt	<= 1'b0;
						state_out	<= IDLE_S;
					end
					else begin
						rdreq_pkt	<= 1'b1;
						state_out	<= READ_FIFO_S;
					end
				end
			endcase	
		end
	end

	
endmodule    
